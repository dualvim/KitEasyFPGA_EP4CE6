module led(output wire [3:0] LED);
	// Acender os 4 LEDs:
	assign LED = 4'b0000;
endmodule
